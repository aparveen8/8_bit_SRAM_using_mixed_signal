* /home/aparveen111/eSim-Workspace/1bitsram/1bitsram.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 08 Oct 2022 10:22:39 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  wl bl Net-_U4-Pad4_ q ayesha_6T_RAM		
U4  Net-_U2-Pad3_ Net-_U2-Pad4_ bl Net-_U4-Pad4_ dac_bridge_2		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ writer_ayesha		
U3  wl din Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
v2  din GND pulse		
v1  wl GND pulse		
SC2  Net-_SC1-Pad1_ q Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__nfet_01v8_lvt		
SC6  dout Net-_SC1-Pad1_ GND GND sky130_fd_pr__nfet_01v8_lvt		
SC3  Net-_SC2-Pad3_ ren GND GND sky130_fd_pr__nfet_01v8_lvt		
v4  ren GND pulse		
v3  Net-_SC1-Pad3_ GND DC		
U6  dout plot_v1		
U5  q plot_v1		
scmode1  SKY130mode		
SC5  dout Net-_SC1-Pad1_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
SC4  Net-_SC1-Pad1_ ren Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		
SC1  Net-_SC1-Pad1_ q Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8_lvt		

.end
